diody zad5
*-------
.LIB EVAL.LIB 

.PARAM RES = 0
*-------
.SUBCKT DZ ZA ZK 

.MODEL DIODE1 D IS=100P N=0.01
.MODEL DIODE2 D IS=100P N=0.01

RZ 2 ZA 20
VZ 1 2 6.7
DZ1 ZK 1 DIODE1
DZ2 ZA ZK DIODE2
.ENDS
*-------	
V1 1 0 10
R1 1 2 500
X1 0 2 DZ
RL 2 0 {RES} 

*-------
.DC V1 6 12 10m
.PROBE
.PLOT DC V(1)
.STEP PARAM RES LIST 1k 2k

.END