zad diody
*-----
.LIB EVAL.LIB
.LIB ANL_MISC.LIB
;D1N750 - zener

*-----
X1 (IN1) 0 (OUT1) 9 (OUT2) XFRM_LIN/CT-SEC

*-----
V1 (IN1) 0 SIN(0 120 60 0 0 0)


D1 (OUT1) 1 D1N4148
D2 0 (OUT2) D1N4148
D3 (OUT2) 1 D1N4148
D4 0 (OUT1) D1N4148

C1 1 0 500u
R1 1 2 200
DZ 0 2 D1N750
RL 2 0 1k

.OP
.TRAN 0 50m 10m


.PROBE
.END
