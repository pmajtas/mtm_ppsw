diody zad3
*-------
.LIB EVAL.LIB 
.PARAM OFFSET =0
.PARAM CAPACITY =0
*-------
V1 1 0 SIN(0 10 1k 0 0 0)
*-------
D1 1 2 D1N4148	
R1 2 0 1k
C1 2 0 {CAPACITY}
*-------

.STEP LIN PARAM CAPACITY 10u 20u 0.2u
.TRAN 0 4m 0.5m 10u
.FOUR 1kHz V(R1)
.PROBE

.END